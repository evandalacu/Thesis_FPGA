module sys_control (

	input clk,
	input en,
	input reset

	)	
	
	
	
endmodule 